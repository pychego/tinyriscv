`timescale 1ns / 1ps

module test ();
    

    reg [3:0] dividend_i;

    initial begin
        dividend_i = -2;
    end


endmodule

